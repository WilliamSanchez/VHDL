library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity SinData is
    port(
        addr : in unsigned(7 downto 0);
        ce : in std_logic;
        out_sin : out unsigned(7 downto 0)
    );
end SinData;

architecture behavioral of SinData is
    type  sin_memory is array (natural range <> ) of unsigned (7 downto 0);
    constant function_sin : sin_memory(0 to 255):=
    ("10000000", "10000011", "10000110", "10001001", "10001100",
     "10001111", "10010010", "10010101", "10011000", "10011100",
     "10011111", "10100010", "10100101", "10101000", "10101011",
     "10101110", "10110000", "10110011", "10110110", "10111001",
     "10111100", "10111111", "11000001", "11000100", "11000111",
     "11001001", "11001100", "11001110", "11010001", "11010011", 
     "11010101", "11011000", "11011010", "11011100", "11011110",
     "11100000", "11100010", "11100100", "11100110", "11101000", 
     "11101010", "11101011", "11101101", "11101111", "11110000",
     "11110010", "11110011", "11110100", "11110110", "11110111",
     "11111000", "11111001", "11111010", "11111011", "11111011", 
     "11111100", "11111101", "11111101", "11111110", "11111110",
     "11111110", "11111111", "11111111", "11111111", "11111111",
     "11111111", "11111111", "11111111", "11111110", "11111110",
     "11111101", "11111101", "11111100", "11111100", "11111011",
     "11111010", "11111001", "11111000", "11110111", "11110110",
     "11110101", "11110100", "11110010", "11110001", "11101111",
     "11101110", "11101100", "11101011", "11101001", "11100111",
     "11100101", "11100011", "11100001", "11011111", "11011101",
     "11011011", "11011001", "11010111", "11010100", "11010010",
     "11001111", "11001101", "11001010", "11001000", "11000101",
     "11000011", "11000000", "10111101", "10111010", "10111000",
     "10110101", "10110010", "10101111", "10101100", "10101001",
     "10100110", "10100011", "10100000", "10011101", "10011010",
     "10010111", "10010100", "10010001", "10001110", "10001010",
     "10000111", "10000100", "10000001", "01111110", "01111011",
     "01111000", "01110101", "01110001", "01101110", "01101011",
     "01101000", "01100101", "01100010", "01011111", "01011100", 
     "01011001", "01010110", "01010011", "01010000", "01001101",
     "01001010", "01000111", "01000101", "01000010", "00111111",
     "00111100", "00111010", "00110111", "00110101", "00110010",
     "00110000", "00101101", "00101011", "00101000", "00100110",
     "00100100", "00100010", "00100000", "00011110", "00011100",
     "00011010", "00011000", "00010110", "00010100", "00010011",
     "00010001", "00010000", "00001110", "00001101", "00001011",
     "00001010", "00001001", "00001000", "00000111", "00000110",
     "00000101", "00000100", "00000011", "00000011", "00000010",
     "00000010", "00000001", "00000001", "00000000", "00000000",
     "00000000", "00000000", "00000000", "00000000", "00000000",
     "00000001", "00000001", "00000001", "00000010", "00000010",
     "00000011", "00000100", "00000100", "00000101", "00000110",
     "00000111", "00001000", "00001001", "00001011", "00001100", 
     "00001101", "00001111", "00010000", "00010010", "00010100",
     "00010101", "00010111", "00011001", "00011011", "00011101",
     "00011111", "00100001", "00100011", "00100101", "00100111",
     "00101010", "00101100", "00101110", "00110001", "00110011",
     "00110110", "00111000", "00111011", "00111110", "00100000",
     "01000011", "01000110", "01001001", "01001100", "01001111",
     "01010001", "01010100", "01010111", "01011010", "01011101",
     "01100000", "01100011", "01100111", "01101010", "01101101",
     "01110000", "01110011", "01110110", "01111001", "01111100",
     "01111100");
    
begin
    out_sin <= function_sin(to_integer(addr)) when ce='0' else (others=>'Z');
end architecture;

--"10000000", "10000011", "10000110", "10001001", "10001100",
--"10001111", "10010010", "10010101", "10011000", "10011100",
--"10011111", "10100010", "10100101", "10101000", "10101011",
--"10101110", "10110000", "10110011", "10110110", "10111001",
--"10111100", "10111111", "11000001", "11000100", "11000111",
--"11001001", "11001100", "11001110", "11010001", "11010011", 
--"11010101", "11011000", "11011010", "11011100", "11011110",
--"11100000", "11100010", "11100100", "11100110", "11101000", 
--"11101010", "11101011", "11101101", "11101111", "11110000",
--"11110010", "11110011", "11110100", "11110110", "11110111",
--"11111000", "11111001", "11111010", "11111011", "11111011", 
--"11111100", "11111101", "11111101", "11111110", "11111110",
--"11111110", "11111111", "11111111", "11111111", "11111111",
--"11111111", "11111111", "11111111", "11111110", "11111110",
--"11111101", "11111101", "11111100", "11111100", "11111011",
--"11111010", "11111001", "11111000", "11110111", "11110110",
--"11110101", "11110100", "11110010", "11110001", "11101111",
--"11101110", "11101100", "11101011", "11101001", "11100111",
--"11100101", "11100011", "11100001", "11011111", "11011101",
--"11011011", "11011001", "11010111", "11010100", "11010010",
--"11001111", "11001101", "11001010", "11001000", "11000101",
--"11000011", "11000000", "10111101", "10111010", "10111000",
--"10110101", "10110010", "10101111", "10101100", "10101001",
--"10100110", "10100011", "10100000", "10011101", "10011010",
--"10010111", "10010100", "10010001", "10001110", "10001010",
--"10000111", "10000100", "10000001", "01111110", "01111011",
--"01111000", "01110101", "01110001", "01101110", "01101011",
--"01101000", "01100101", "01100010", "01011111", "01011100", 
--"01011001", "01010110", "01010011", "01010000", "01001101",
--"01001010", "01000111", "01000101", "01000010", "00111111",
--"00111100", "00111010", "00110111", "00110101", "00110010",
--"00110000", "00101101", "00101011", "00101000", "00100110",
--"00100100", "00100010", "00100000", "00011110", "00011100",
--"00011010", "00011000", "00010110", "00010100", "00010011",
--"00010001", "00010000", "00001110", "00001101", "00001011",
--"00001010", "00001001", "00001000", "00000111", "00000110",
--"00000101", "00000100", "00000011", "00000011", "00000010",
--"00000010", "00000001", "00000001", "00000000", "00000000",
--"00000000", "00000000", "00000000", "00000000", "00000000",
--"00000001", "00000001", "00000001", "00000010", "00000010",
--"00000011", "00000100", "00000100", "00000101", "00000110",
--"00000111", "00001000", "00001001", "00001011", "00001100", 
--"00001101", "00001111", "00010000", "00010010", "00010100",
--"00010101", "00010111", "00011001", "00011011", "00011101",
--"00011111", "00100001", "00100011", "00100101", "00100111",
--"00101010", "00101100", "00101110", "00110001", "00110011",
--"00110110", "00111000", "00111011", "00111110", "00100000",
--"01000011", "01000110", "01001001", "01001100", "01001111",
--"01010001", "01010100", "01010111", "01011010", "01011101",
--"01100000", "01100011", "01100111", "01101010", "01101101",
--"01110000", "01110011", "01110110", "01111001", "01111100",
